library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity laelaps_four_legs_duplicate_ip_v1_0 is
	generic (  --This is the top module of our IP and hence the values defined here are the ones that determine the rest of the generic variables in all subcomponents
		-- Users to add parameters here
        sys_clk : INTEGER := 90_909_088;            --system clock frequency in Hz
        pwm_frequency   : INTEGER := 20_000;        --PWM switching frequency in Hz
        bits_resolution : INTEGER := 14;            --bits of resolution setting the duty cycle
        phases          : INTEGER := 1; 
        bits            : INTEGER := 18;            --number of bits for encoder's counts
        hip_ratio_numerator   : INTEGER := 1029;    --numerator of the gear ratio of the Hip motor-gearhead
        hip_ratio_divisor : INTEGER := 13;          --divisor of the gear ratio of the Hip motor-gearhead
        knee_ratio_numerator : INTEGER := 98;       --numerator of the gear ratio of the Knee motor-gearhead
        knee_ratio_divisor : INTEGER := 1;          --divisor of the gear ratio of the Hip motor-gearhead
		-- User parameters ends
		-- Do not modify the parameters beyond this line


		-- Parameters of Axi Slave Bus Interface S00_AXI
		C_S00_AXI_DATA_WIDTH	: integer	:= 32;
		C_S00_AXI_ADDR_WIDTH	: integer	:= 7
	);
	port (
		-- Users to add ports here
        jb_p0 : in std_logic;   --A1 of first leg                      
        jb_n0 : in std_logic;   --B1 of first leg
        jb_p1 : in std_logic;   --A2 of first leg
        jb_n1 : in std_logic;   --B2 of first leg
        jb_p2 : out std_logic;  --DIR1 of first leg
        jb_n2 : out std_logic;  --PWM1 of first leg
        jb_p3 : out std_logic;  --DIR2 of first leg
        jb_n3 : out std_logic;  --PWM2 of first leg
        
        jc_p0 : in std_logic;   --A1 of second leg                       
        jc_n0 : in std_logic;   --B1 of second leg
        jc_p1 : in std_logic;   --A2 of second leg
        jc_n1 : in std_logic;   --B2 of second leg
        jc_p2 : out std_logic;  --DIR1 of second leg
        jc_n2 : out std_logic;  --PWM1 of second leg
        jc_p3 : out std_logic;  --DIR2 of second leg
        jc_n3 : out std_logic;  --PWM2 of second leg
        
        jd_p0 : in std_logic;   --A1 of third leg                      
        jd_n0 : in std_logic;   --B1 of third leg
        jd_p1 : in std_logic;   --A2 of third leg
        jd_n1 : in std_logic;   --B2 of third leg
        jd_p2 : out std_logic;  --DIR1 of third leg
        jd_n2 : out std_logic;  --PWM1 of third leg
        jd_p3 : out std_logic;  --DIR2 of third leg
        jd_n3 : out std_logic;  --PWM2 of third leg
        
        je_p0 : in std_logic;   --A1 of fourth leg                       
        je_n0 : in std_logic;   --B1 of fourth leg
        je_p1 : in std_logic;   --A2 of fourth leg
        je_n1 : in std_logic;   --B2 of fourth leg
        je_p2 : out std_logic;  --DIR1 of fourth leg
        je_n2 : out std_logic;  --PWM1 of fourth leg
        je_p3 : out std_logic;  --DIR2 of fourth leg
        je_n3 : out std_logic;  --PWM2 of fourth leg
        led : out std_logic_vector(3 downto 0);     --leds of Zybo Board
        sw : in std_logic_vector(3 downto 0);       --switches of Zybo Board
		-- User ports ends
		-- Do not modify the ports beyond this line


		-- Ports of Axi Slave Bus Interface S00_AXI
		s00_axi_aclk	: in std_logic;
		s00_axi_aresetn	: in std_logic;
		s00_axi_awaddr	: in std_logic_vector(C_S00_AXI_ADDR_WIDTH-1 downto 0);
		s00_axi_awprot	: in std_logic_vector(2 downto 0);
		s00_axi_awvalid	: in std_logic;
		s00_axi_awready	: out std_logic;
		s00_axi_wdata	: in std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
		s00_axi_wstrb	: in std_logic_vector((C_S00_AXI_DATA_WIDTH/8)-1 downto 0);
		s00_axi_wvalid	: in std_logic;
		s00_axi_wready	: out std_logic;
		s00_axi_bresp	: out std_logic_vector(1 downto 0);
		s00_axi_bvalid	: out std_logic;
		s00_axi_bready	: in std_logic;
		s00_axi_araddr	: in std_logic_vector(C_S00_AXI_ADDR_WIDTH-1 downto 0);
		s00_axi_arprot	: in std_logic_vector(2 downto 0);
		s00_axi_arvalid	: in std_logic;
		s00_axi_arready	: out std_logic;
		s00_axi_rdata	: out std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
		s00_axi_rresp	: out std_logic_vector(1 downto 0);
		s00_axi_rvalid	: out std_logic;
		s00_axi_rready	: in std_logic
	);
end laelaps_four_legs_duplicate_ip_v1_0;

architecture arch_imp of laelaps_four_legs_duplicate_ip_v1_0 is

	-- component declaration
	component laelaps_four_legs_duplicate_ip_v1_0_S00_AXI is
		generic (
        sys_clk         : INTEGER := 100_000_000;       --system clock frequency in Hz
        pwm_frequency   : INTEGER := 20_000;            --PWM switching frequency in Hz
        bits_resolution : INTEGER := 14;                --bits of resolution setting the duty cycle
        phases          : INTEGER := 1; 
        bits            : INTEGER := 18;                --number of bits for encoder's counts
        hip_ratio_numerator   : INTEGER := 1029;    --numerator of the gear ratio of the Hip motor-gearhead
        hip_ratio_divisor : INTEGER := 13;          --divisor of the gear ratio of the Hip motor-gearhead
        knee_ratio_numerator : INTEGER := 98;      --numerator of the gear ratio of the Knee motor-gearhead
        knee_ratio_divisor : INTEGER := 1;          --divisor of the gear ratio of the Hip motor-gearhead
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		C_S_AXI_ADDR_WIDTH	: integer	:= 7
		);
		port (
        jb_p0 : in std_logic;   --A1 of first leg                      
        jb_n0 : in std_logic;   --B1 of first leg
        jb_p1 : in std_logic;   --A2 of first leg
        jb_n1 : in std_logic;   --B2 of first leg
        jb_p2 : out std_logic;  --DIR1 of first leg
        jb_n2 : out std_logic;  --PWM1 of first leg
        jb_p3 : out std_logic;  --DIR2 of first leg
        jb_n3 : out std_logic;  --PWM2 of first leg
        jc_p0 : in std_logic;   --A1 of second leg                       
        jc_n0 : in std_logic;   --B1 of second leg
        jc_p1 : in std_logic;   --A2 of second leg
        jc_n1 : in std_logic;   --B2 of second leg
        jc_p2 : out std_logic;  --DIR1 of second leg
        jc_n2 : out std_logic;  --PWM1 of second leg
        jc_p3 : out std_logic;  --DIR2 of second leg
        jc_n3 : out std_logic;  --PWM2 of second leg
        jd_p0 : in std_logic;   --A1 of third leg                      
        jd_n0 : in std_logic;   --B1 of third leg
        jd_p1 : in std_logic;   --A2 of third leg
        jd_n1 : in std_logic;   --B2 of third leg
        jd_p2 : out std_logic;  --DIR1 of third leg
        jd_n2 : out std_logic;  --PWM1 of third leg
        jd_p3 : out std_logic;  --DIR2 of third leg
        jd_n3 : out std_logic;  --PWM2 of third leg
        je_p0 : in std_logic;   --A1 of fourth leg                       
        je_n0 : in std_logic;   --B1 of fourth leg
        je_p1 : in std_logic;   --A2 of fourth leg
        je_n1 : in std_logic;   --B2 of fourth leg
        je_p2 : out std_logic;  --DIR1 of fourth leg
        je_n2 : out std_logic;  --PWM1 of fourth leg
        je_p3 : out std_logic;  --DIR2 of fourth leg
        je_n3 : out std_logic;  --PWM2 of fourth leg
        led : out std_logic_vector(3 downto 0);
        sw : in std_logic_vector(3 downto 0);
		S_AXI_ACLK	: in std_logic;
		S_AXI_ARESETN	: in std_logic;
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		S_AXI_AWVALID	: in std_logic;
		S_AXI_AWREADY	: out std_logic;
		S_AXI_WDATA	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_WSTRB	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		S_AXI_WVALID	: in std_logic;
		S_AXI_WREADY	: out std_logic;
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		S_AXI_BVALID	: out std_logic;
		S_AXI_BREADY	: in std_logic;
		S_AXI_ARADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		S_AXI_ARVALID	: in std_logic;
		S_AXI_ARREADY	: out std_logic;
		S_AXI_RDATA	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		S_AXI_RVALID	: out std_logic;
		S_AXI_RREADY	: in std_logic
		);
	end component laelaps_four_legs_duplicate_ip_v1_0_S00_AXI;

begin

-- Instantiation of Axi Bus Interface S00_AXI
laelaps_four_legs_duplicate_ip_v1_0_S00_AXI_inst : laelaps_four_legs_duplicate_ip_v1_0_S00_AXI
	generic map (
        sys_clk => sys_clk,                      --system clock frequency in Hz
        pwm_frequency   => pwm_frequency,       --PWM switching frequency in Hz
        bits_resolution => bits_resolution,     --bits of resolution setting the duty cycle
        phases    => phases, 
        bits => bits,
        hip_ratio_numerator => hip_ratio_numerator,
        hip_ratio_divisor => hip_ratio_divisor,
        knee_ratio_numerator => knee_ratio_numerator,
        knee_ratio_divisor => knee_ratio_divisor,
		C_S_AXI_DATA_WIDTH	=> C_S00_AXI_DATA_WIDTH,
		C_S_AXI_ADDR_WIDTH	=> C_S00_AXI_ADDR_WIDTH
	)
	port map (
        jb_p0 => jb_p0,
        jb_n0 => jb_n0,
        jb_p1 => jb_p1,
        jb_n1 => jb_n1,
        jb_p2 => jb_p2,
        jb_n2 => jb_n2,
        jb_n3 => jb_n3,
        jb_p3 => jb_p3,
        jc_p0 => jc_p0,
        jc_n0 => jc_n0,
        jc_p1 => jc_p1,
        jc_n1 => jc_n1,
        jc_p2 => jc_p2,
        jc_n2 => jc_n2,
        jc_n3 => jc_n3,
        jc_p3 => jc_p3,
        jd_p0 => jd_p0,
        jd_n0 => jd_n0,
        jd_p1 => jd_p1,
        jd_n1 => jd_n1,
        jd_p2 => jd_p2,
        jd_n2 => jd_n2,
        jd_n3 => jd_n3,
        jd_p3 => jd_p3,
        je_p0 => je_p0,
        je_n0 => je_n0,
        je_p1 => je_p1,
        je_n1 => je_n1,
        je_p2 => je_p2,
        je_n2 => je_n2,
        je_n3 => je_n3,
        je_p3 => je_p3,
        led => led,
        sw => sw,
		S_AXI_ACLK	=> s00_axi_aclk,
		S_AXI_ARESETN	=> s00_axi_aresetn,
		S_AXI_AWADDR	=> s00_axi_awaddr,
		S_AXI_AWPROT	=> s00_axi_awprot,
		S_AXI_AWVALID	=> s00_axi_awvalid,
		S_AXI_AWREADY	=> s00_axi_awready,
		S_AXI_WDATA	=> s00_axi_wdata,
		S_AXI_WSTRB	=> s00_axi_wstrb,
		S_AXI_WVALID	=> s00_axi_wvalid,
		S_AXI_WREADY	=> s00_axi_wready,
		S_AXI_BRESP	=> s00_axi_bresp,
		S_AXI_BVALID	=> s00_axi_bvalid,
		S_AXI_BREADY	=> s00_axi_bready,
		S_AXI_ARADDR	=> s00_axi_araddr,
		S_AXI_ARPROT	=> s00_axi_arprot,
		S_AXI_ARVALID	=> s00_axi_arvalid,
		S_AXI_ARREADY	=> s00_axi_arready,
		S_AXI_RDATA	=> s00_axi_rdata,
		S_AXI_RRESP	=> s00_axi_rresp,
		S_AXI_RVALID	=> s00_axi_rvalid,
		S_AXI_RREADY	=> s00_axi_rready
	);

	-- Add user logic here

	-- User logic ends

end arch_imp;

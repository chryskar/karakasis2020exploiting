----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/20/2018 03:50:34 PM
-- Design Name: 
-- Module Name: qei - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity qei is
    generic(
            sys_clk         : INTEGER := 100_000_000;           --system clock frequency in Hz
            bits            : INTEGER := 18;                    --number of ratio bits
            ratio_numerator : INTEGER := 98;                    --numerator of the gear ratio of the motor-gearhead
            ratio_divisor   : INTEGER := 1                      --divisor of the gear ratio of the motor-gearhead
            ); 
    Port ( 
           QEA : in STD_LOGIC;                                  --The A signal as generated from the encoder
           Index : in STD_LOGIC;                                --The Index signal as generated from the encoder
           QEB : in STD_LOGIC;                                  --The B signal as generated from the encoder
           Clk : in STD_LOGIC;                                  --The Clock Signal
           Count_out : out STD_LOGIC_VECTOR (bits-1 downto 0);  --The Calculated Position of the Motor in Counts
           vel_sign : out STD_LOGIC;                            --The Calculated Sign of the Motor's Velocity
           velocity : out STD_LOGIC_VECTOR  (31 downto 0)       --The Calculated Value of the Motor's Velocity
           );
end qei;

architecture Behavioral of qei is
signal F1_out : STD_LOGIC;
signal F2_out : STD_LOGIC;
signal F3_out : STD_LOGIC;
signal c_clk : STD_LOGIC;
signal r_clk : STD_LOGIC;
signal clk2 : STD_LOGIC:= '0';
signal r_count : STD_LOGIC;
signal temp_count : STD_LOGIC_VECTOR (bits-1 downto 0);
signal temp_dir : std_logic;

COMPONENT filter IS                                             --Declaration of the "filter" Component
  PORT(
		QEX : in STD_LOGIC;                                     -- First input is a 1-bit signal generated from an encoder, either the A,B or Index
        clk : in STD_LOGIC;                                     -- For synchronization reasons a 1-bit clock signal is linked
        fout : out STD_LOGIC                                    -- The output of our system is a 1-bit signal
		);
END COMPONENT;

COMPONENT encoder IS                                            --Declaration of the "encoder" Component
    generic(            --The actual values of the generic variables are specified in Line 141-145
        bits  : INTEGER := 18;                                  --number of ratio bits
        ratio_numerator : INTEGER := 98;                        --numerator of the gear ratio of the motor-gearhead
        ratio_divisor : INTEGER := 1                            --divisor of the gear ratio of the motor-gearhead
        ); 
  PORT(
        QuadA : in STD_LOGIC;                                   --Filtered 1-Bit Signal A from the encoder
        QuadB : in STD_LOGIC;                                   --Filtered 1-Bit Signal B from the encoder
        Index : in STD_LOGIC;                                   --Filtered 1-Bit Signal Index from the encoder
        Clk : in STD_LOGIC;                                     --1-Bit Clock Signal for synchronization reasons
        DIR : out STD_LOGIC;                                    --Output 1-Bit Signal that shows the direction of motion (Clockwise or Anti-Clockwise)
        Position : out STD_LOGIC_VECTOR (bits-1 downto 0)       --Output bits-Bits Signal that shows the position of the motor in counts
		);
END COMPONENT;

COMPONENT vel_qei IS
    generic(            --The actual values of the generic variables are specified in Line 156-160
    sys_clk         : INTEGER := 100_000_000;                   --system clock frequency in Hz
    bits            : INTEGER := 18;                            --number of ratio bit
    ratio_numerator : INTEGER := 98;                            --numerator of the gear ratio of the motor-gearhead
    ratio_divisor   : INTEGER := 1                              --divisor of the gear ratio of the motor-gearhead
    ); 
  Port (   DIR_in : in STD_LOGIC;                               --Direction of Motion
           count_in : in STD_LOGIC_VECTOR (bits-1 downto 0);    --Position of Motor
           Clk : in STD_LOGIC;                                  --Clock Signal
           velocity_sign : out std_logic;                       --The sign of the estimated motor's velocity
           velocity_temp : out std_logic_vector (31 downto 0)); --The motor's estimated velocity
END COMPONENT;

begin

p_200_kHZ : process (Clk) is                                    --This process creates a four times slower clock signal than the Clk Signal 
  begin
    if rising_edge(Clk) then                                    --Everytime the Clk signal changes from '0' to '1'
      if r_count = '1' then                                     --Counter of changes in the Clk Signal
        clk2 <= not clk2;                                       --The slow clock signal changes every second time a rising edge occurs in the fast clock
        r_count    <= '0';                                      --Update of the Counter of changes in the Clk Signal
      else
        r_count <= '1';                                         --Update of the Counter of changes in the Clk Signal
      end if;
    end if;
  end process p_200_kHZ;
  
F1: filter                                                      --Utilization of the first "filter" component for the A signal of the encoder
PORT MAP 
(
QEX  => QEA,                                                    --The A signal of the encoder is supplied to the filter block
clk  => Clk,                                                    --The fast clock is supplied to the filter block
fout => F1_out                                                  --The filter blocks outputs the stable and filtered A signal
);

F2: filter                                                      --Utilization of the second "filter" component for the B signal of the encoder
PORT MAP   
(
QEX  => QEB,                                                    --The B signal of the encoder is supplied to the filter block
clk  => Clk,                                                    --The fast clock is supplied to the filter block
fout => F2_out                                                  --The filter blocks outputs the stable and filtered B signal
);

F3: filter                                                      --Utilization of the third "filter" component for the Index signal of the encoder  
PORT MAP 
(
QEX  => Index,                                                  --The Index signal of the encoder is supplied to the filter block
clk  => Clk,                                                    --The fast clock is supplied to the filter block
fout => F3_out                                                  --The filter blocks outputs the stable and filtered Index signal
);

E1: encoder                                                     --Utilization of the "encoder" component for the calculation of the Motor's Position
generic map (                                                   --Generic Variables are defined here according to the values of the signals on the right 
bits => bits,                                                   --which will be specified when the "qei" block will be called as 
ratio_numerator => ratio_numerator,                             --a component by another function. Otherwise, they will be equal to the top definition (See Line 36-41)
ratio_divisor => ratio_divisor) 
PORT MAP 
(
QuadA  => F1_out,                                               --The filtered signal A is given as input to the "encoder" component
QuadB  => F2_out,                                               --The filtered signal B is given as input to the "encoder" component
Index => F3_out,                                                --The filtered signal Index is given as input to the "encoder" component
    Clk  => clk2,                                                   --The slow clock is supplied to the "encoder" block
DIR => temp_dir,                                                --The "encoder" block outputs the Motion's Direction
Position => temp_count                                          --The "encoder" block outputs the Motor's Position in counts
);

V1: vel_qei                                                     --Utilization of the "vel_qei" component for the calculation of the Motor's Velocity
generic map (                                                   --Generic Variables are defined here according to the values of the signals on the right 
sys_clk => sys_clk,                                             --which will be specified when the "qei" block will be called as 
bits => bits, --number of ratio bit                             --a component by another function. Otherwise, they will be equal to the top definition (See Line 36-41)
ratio_numerator => ratio_numerator,
ratio_divisor => ratio_divisor
)
PORT MAP 
(
DIR_in => temp_dir,                                             --The calculated Motion's Direction is given as input to the "vel_qei" component
count_in => temp_count,                                         --The calculated Motor's Position is given as input to the "vel_qei" component
Clk => clk2,                                                    --The slow clock is supplied to the "vel_qei" block
velocity_sign => vel_sign,                                      --The "vel_qei" block outputs the velocity's sign as one of the "qei" block's outputs
velocity_temp => velocity                                       --The "vel_qei" block outputs the velocity's value as one of the "qei" block's outputs
);

Count_out <= temp_count;                                        --The "qei" block outputs the Motor's Position
end Behavioral;

----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/19/2018 07:00:56 PM
-- Design Name: 
-- Module Name: filter - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

--This block receives as inputs the signals generated from the encoders and checks whether they are stable or not. 
--If yes, then they are transferred to the next processing level. Otherwise, the output is not modified.

entity filter is
    Port ( QEX : in STD_LOGIC;                                  -- First input is a 1-bit signal generated from an encoder, either the A,B or Index
           clk : in STD_LOGIC;                                  -- For synchronization reasons a 1-bit clock signal is linked
           fout : out STD_LOGIC);                               -- The output of our system is a 1-bit signal
end filter;

architecture Behavioral of filter is

signal QEX_Delayed: STD_LOGIC_VECTOR(2 downto 0) := "000";      -- A 3-bit auxiliary signal

begin
process (clk)                                                   -- Everytime the "clk" changes, the code inside the process is executed
begin
    if (clk='1' and clk'event) then                             -- This check is for the detection of a rising edge in the clock signal
        QEX_Delayed <= (QEX_Delayed(1), QEX_Delayed(0), QEX);   -- Store the new QEX input in the first bit of the QEX_Delayed signal, while shifting the previous first and second bits to the current third and second
        if QEX_Delayed = "000" then                             -- If the last three samples of the input are equal to each other and to zero, the signal is considered stable and the output is set to zero
            fout <= '0';
        elsif QEX_Delayed = "111" then                          -- If the last three samples of the input are equal to each other and to one, the signal is considered stable and the output is set to one
            fout <= '1';
        end if;
    end if;
end process;

end Behavioral;

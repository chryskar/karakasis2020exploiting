----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07/30/2018 02:08:24 PM
-- Design Name: 
-- Module Name: vel_qei - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use IEEE.std_logic_arith.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
    
entity vel_qei is
    generic(            --The actual values of the generic variables are not the following (18,98 and 1) but they will be specified by the module that utilizes the encoder code as a component (See "qei.vhd")
        sys_clk         : INTEGER := 100_000_000;                       --system clock frequency in Hz
        bits            : INTEGER := 18;                                --number of ratio bit
        ratio_numerator : INTEGER := 98;                                --numerator of the gear ratio of the motor-gearhead
        ratio_divisor   : INTEGER := 1                                  --divisor of the gear ratio of the motor-gearhead
        );     
    Port ( DIR_in : in STD_LOGIC;                                       --Direction of Motion
           count_in : in STD_LOGIC_VECTOR (bits-1 downto 0);            --Position of Motor
           Clk : in STD_LOGIC;                                          --Clock Signal
           velocity_sign : out std_logic;                               --The sign of the estimated motor's velocity
           velocity_temp : out std_logic_vector (31 downto 0));         --The motor's estimated velocity
end vel_qei;

architecture Behavioral of vel_qei is
CONSTANT  vel_constant  :  INTEGER :=  31415927;                        --First constant of the Velocity Estimation Equation
CONSTANT  f_FPGA  :  INTEGER :=  sys_clk/1000000;                       --Second constant of the Velocity Estimation Equation
CONSTANT  temp1 :  INTEGER := vel_constant*ratio_divisor/ratio_numerator;   --Third constant of the Velocity Estimation Equation
CONSTANT  vel_numerator  :  INTEGER :=  temp1*f_fpga;                   --Fourth constant of the Velocity Estimation Equation
CONSTANT  zero_constant  :  INTEGER :=  vel_numerator/10;               --Fifth constant of the Velocity Estimation Equation
signal sum_QCLK: STD_LOGIC_VECTOR(2 downto 0) := (others => '0');
signal DT : STD_LOGIC_VECTOR (31 downto 0) := std_logic_vector(to_unsigned(vel_numerator,32));   --max value of DT in binary
signal error_flag : std_logic := '0';                                               --Initialization
signal DIR_change : std_logic := '0';                                               --Initialization
signal temp_DIR : std_logic := '1';                                                 --Initialization
signal A_trunc : STD_LOGIC_VECTOR (31 downto 0):= (others => '0');                  --Initialization
signal B_trunc : STD_LOGIC_VECTOR (31 downto 0):= (others => '1');                  --Initialization
signal DIR_temp : std_logic:='1';                                                   --Initialization
signal vel_flag : std_logic_vector(1 downto 0):="00";                               --Initialization
signal count_last : STD_LOGIC_VECTOR (bits-1 downto 0):=(others => '0');            --Initialization

begin
process (Clk)                                                           --Everytime a change occurs in the Clock signal the code inside the process are being executed
begin
    if Clk='1' and Clk'event then                                       --Rising Edge Detection of the Clock Signal
        DT <= DT + 1;                                                   --Counter of the Clock Cycles
        if DT = std_logic_vector(to_unsigned(zero_constant,DT'length)) then --When the Clock Cycles Counter reaches this value, the velocity is practically zero
            error_flag <= '1';                                          --This informs us that later on we should set the velocity to zero
        end if;
        if DIR_in /= DIR_temp then                                      --Change in direction, DIR_temp holds the previous clock value of the DIR signal
            DIR_temp <= DIR_in;                                         --Update of the Direction Signal for comparison with the next one (It takes a cycle to see the new value)
            if DIR_in /= temp_DIR then                                  --Comparion with current direction
                DIR_change <= '1';                                      --Flag signal to notify the change of direction
            end if;
        end if;
        if (count_in /= count_last) then                                --Change in the Motor's Position
            count_last <= count_in;                                     --Update of the temp signal that keeps track of the Position
            if sum_QCLK < "011" then                                    --Chech whether 4 changes have occured in the Position Signal
                sum_QCLK <= sum_QCLK + 1;                               --If not, increase of the changes counter
            else                                                        --Otherwise, we check for overflow
                if error_flag = '1' then                                --Check whether the velocity should be set to zero
                    B_trunc(31 downto 0) <= (others => '1');            --By setting the Divisor to maximum the velocity will become zero
                    error_flag <= '0';                                  --Clear the overflow error flag
                else                                                    --No overflow
                    B_trunc(31 downto 0) <= DT;                         --Updating the Divisor with the counted Clock Cycles that occured between the four changes in the Position Signal
                end if;
                                                                        --Check for change in direction
                if DIR_change = '1' then                                --change of direction
                    vel_flag <= "00";                                   --Flag signal for command in Line 115 to set Velocity to zero
                    DIR_change <= '0';                                  --Clear direction flag
                    temp_DIR <= DIR_in;                                 --Update of the Direction output signals (See Line 120)
                else                                                    --no change in direction 
                                                                        --velocity <= count/DT; 
                    if DT = "00000000000000000000000000000000" then     --check if devisor is equal to zero.
                        B_trunc(31 downto 0) <= (others => '1');        --velocity = 0
                        vel_flag <= "01";                               --Flag signal for command in Line 115 to set Velocity to Maximum
                    else                                                --if not, complete the division
                        A_trunc(31 downto 0) <= std_logic_vector(to_unsigned(vel_numerator,A_trunc'length)); --Update the dividend
                        vel_flag <= "10";                               --Flag signal for command in Line 115 to execute the division and calculate the Velocity
                    end if;
                end if;
                sum_QCLK <= (others => '0');                            --Clear the counter that keeps track of the Position Signal's changes
                DT <= (others => '0');                                  --Clear the Clock Cycles Counter
            end if;
        end if;
    end if;    
end process;

velocity_temp <= std_logic_vector ( unsigned(A_trunc) / unsigned(B_trunc) ) when vel_flag="10" and error_flag = '0' else
                  (others => '0') when vel_flag="00" or error_flag = '1' else
                  (others => '1');                        --In the first case, the division is completed and the velocity is estimated
                                                          --In the second case, the velocity is set to zero
                                                          --In the third case, the velocity is set to Maximum Value
velocity_sign <= temp_DIR;                                --The two signals are always equal to each other
end Behavioral;

----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/14/2018 03:41:20 PM
-- Design Name: 
-- Module Name: encoder - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity encoder is
    generic(                                --The actual values of the generic variables are not the following (18,98 and 1) but they will be specified by the module that utilizes the encoder code as a component (See "qei.vhd")
    bits  : INTEGER := 18;                  --number of ratio bits 
    ratio_numerator : INTEGER := 98;        --numerator of the gear ratio of the motor-gearhead
    ratio_divisor : INTEGER := 1            --divisor of the gear ratio of the motor-gearhead
    ); 
    Port ( 
           QuadA : in STD_LOGIC;            --Filtered 1-Bit Signal A from the encoder
           QuadB : in STD_LOGIC;            --Filtered 1-Bit Signal B from the encoder
           Index : in STD_LOGIC;            --Filtered 1-Bit Signal Index from the encoder
           Clk : in STD_LOGIC;              --1-Bit Clock Signal for synchronization reasons
           DIR : out STD_LOGIC;             --Output 1-Bit Signal that shows the direction of motion (Clockwise or Anti-Clockwise)
           Position : out STD_LOGIC_VECTOR (bits-1 downto 0) --Output bits-Bits Signal that shows the position of the motor in counts
    );
end encoder;

architecture Behavioral of encoder is
CONSTANT  max_value     :  INTEGER := ratio_numerator*2000/ratio_divisor;   --Auxiliary Constant of the maximum value that a Position signal can reach 
signal QuadA_Delayed: STD_LOGIC_VECTOR(2 downto 0) := "000";                --Auxiliary 3-bit Signal that stores the last three values of the A input
signal QuadB_Delayed: STD_LOGIC_VECTOR(2 downto 0) := "000";                --Auxiliary 3-bit Signal that stores the last three values of the B input
 
signal Count_Enable_temp: STD_LOGIC;                                        --Auxiliary Intermediate 1-bit Signal
signal Count_Direction_temp: STD_LOGIC;                                     --Auxiliary Intermediate 1-bit Signal
 
signal Count: STD_LOGIC_VECTOR(bits-1 downto 0) := (others => '0');         --Intermediate Signal for the Position Signal
begin
 
process (Clk,Index)                                                             --The code inside the Process will be executed everytime a chance occurs in either the Clock or Index Signals
begin
    if Index='1' then                                                               --If the Index Signal is equal to 1, the counter has to reset to zero.
        Count <= (others => '0' );                                                  --The Count Signal is used as a substitute for the Position Signal (See lines 72 and 89) 
	elsif Clk='1' and Clk'event then                                                --Rising Edge Detection of the Clock Signal
		QuadA_Delayed <= (QuadA_Delayed(1), QuadA_Delayed(0), QuadA);               --Storing and Update of the Last three samples of the A input     
		QuadB_Delayed <= (QuadB_Delayed(1), QuadB_Delayed(0), QuadB);               --Storing and Update of the last three samples of the B input
        if Count_Enable_temp='1' then                                               --Check whether the Inputs have changed during the last two samples (For the Definition of the Count_Enable_temp see Line 90)
            if Count_Direction_temp='1' then                                        --If Direction is Positive, we increase the counter (See Line 92)
                if Count < max_value then                                           --Check whether the Signal has reached maximum value
                    Count <= Count + 1;                                             --If not, the Count increases (We could not use the Position Signal instead of the Count, due to the fact that a Signal declared as Output cannot be used as an input to a command)
                    DIR <= '1';                                                     --and the Direction Signal is set to 1 and states Positive Motion
                else                                                                --If yes, the Count resets to zero
                    Count <= (others => '0' ); 
                end if;
            else                                                                    --If Direction is Negative, we decrease the counter (See Line 92)
                if Count > 0 then                                                   --Check whether the Signal has reached minimum value 
                    Count <= Count - 1;                                             --If not, the Count decreases (We could not use the Position Signal instead of the Count, due to the fact that a Signal declared as Output cannot be used as an input to a command)
                    DIR <= '0';                                                     --and the Direction Signal is set to 0 and states Negative Motion
                else 
                    Count <= std_logic_vector(to_unsigned(max_value,Count'length)); --If yes, the Count resets to the maximum value
                end if;
            end if;
        end if;
	end if;
end process;
                                                                                    --All commands outside the process field are being executed constantly
Position <= Count;                                                                  --Constantly the Position signal is equal to the Count signal
Count_Enable_temp <= QuadA_Delayed(1) xor QuadA_Delayed(2) xor QuadB_Delayed(1)
				xor QuadB_Delayed(2);                                           --If both Inputs have not changed during the last two samples, the system's output remains the same and hence there is no reason for computation
Count_Direction_temp <= QuadA_Delayed(1) xor QuadB_Delayed(2);                  --According to this signal we can deduce the direction of motion for the motor
end Behavioral;

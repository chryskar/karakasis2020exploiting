library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

    entity laelaps_four_legs_duplicate_ip_v1_0_S00_AXI is
	generic (
		-- Users to add parameters here
        sys_clk         : INTEGER := 100_000_000;   --system clock frequency in Hz
        pwm_frequency   : INTEGER := 20_000;        --PWM switching frequency in Hz
        bits_resolution : INTEGER := 14;            --bits of resolution setting the duty cycle
        phases          : INTEGER := 1; 
        bits            : INTEGER := 18;            --number of bits for encoder's counts
        hip_ratio_numerator   : INTEGER := 1029;    --numerator of the gear ratio of the Hip motor-gearhead
        hip_ratio_divisor : INTEGER := 13;          --divisor of the gear ratio of the Hip motor-gearhead
        knee_ratio_numerator : INTEGER := 98;       --numerator of the gear ratio of the Knee motor-gearhead
        knee_ratio_divisor : INTEGER := 1;          --divisor of the gear ratio of the Hip motor-gearhead
		-- User parameters ends
		-- Do not modify the parameters beyond this line

		-- Width of S_AXI data bus
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		-- Width of S_AXI address bus
		C_S_AXI_ADDR_WIDTH	: integer	:= 7
	);
	port (
		-- Users to add ports here
        jb_p0 : in std_logic;   --A1 of first leg                      
        jb_n0 : in std_logic;   --B1 of first leg
        jb_p1 : in std_logic;   --A2 of first leg
        jb_n1 : in std_logic;   --B2 of first leg
        jb_p2 : out std_logic;  --DIR1 of first leg
        jb_n2 : out std_logic;  --PWM1 of first leg
        jb_p3 : out std_logic;  --DIR2 of first leg
        jb_n3 : out std_logic;  --PWM2 of first leg
        
        jc_p0 : in std_logic;   --A1 of second leg                       
        jc_n0 : in std_logic;   --B1 of second leg
        jc_p1 : in std_logic;   --A2 of second leg
        jc_n1 : in std_logic;   --B2 of second leg
        jc_p2 : out std_logic;  --DIR1 of second leg
        jc_n2 : out std_logic;  --PWM1 of second leg
        jc_p3 : out std_logic;  --DIR2 of second leg
        jc_n3 : out std_logic;  --PWM2 of second leg
        
        jd_p0 : in std_logic;   --A1 of third leg                      
        jd_n0 : in std_logic;   --B1 of third leg
        jd_p1 : in std_logic;   --A2 of third leg
        jd_n1 : in std_logic;   --B2 of third leg
        jd_p2 : out std_logic;  --DIR1 of third leg
        jd_n2 : out std_logic;  --PWM1 of third leg
        jd_p3 : out std_logic;  --DIR2 of third leg
        jd_n3 : out std_logic;  --PWM2 of third leg
        
        je_p0 : in std_logic;   --A1 of fourth leg                       
        je_n0 : in std_logic;   --B1 of fourth leg
        je_p1 : in std_logic;   --A2 of fourth leg
        je_n1 : in std_logic;   --B2 of fourth leg
        je_p2 : out std_logic;  --DIR1 of fourth leg
        je_n2 : out std_logic;  --PWM1 of fourth leg
        je_p3 : out std_logic;  --DIR2 of fourth leg
        je_n3 : out std_logic;  --PWM2 of fourth leg
        led : out std_logic_vector(3 downto 0);     --leds of Zybo Board
        sw : in std_logic_vector(3 downto 0);       --switches of Zybo Board
		-- User ports ends
		-- Do not modify the ports beyond this line

		-- Global Clock Signal
		S_AXI_ACLK	: in std_logic;
		-- Global Reset Signal. This Signal is Active LOW
		S_AXI_ARESETN	: in std_logic;
		-- Write address (issued by master, acceped by Slave)
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		-- Write channel Protection type. This signal indicates the
    		-- privilege and security level of the transaction, and whether
    		-- the transaction is a data access or an instruction access.
		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		-- Write address valid. This signal indicates that the master signaling
    		-- valid write address and control information.
		S_AXI_AWVALID	: in std_logic;
		-- Write address ready. This signal indicates that the slave is ready
    		-- to accept an address and associated control signals.
		S_AXI_AWREADY	: out std_logic;
		-- Write data (issued by master, acceped by Slave) 
		S_AXI_WDATA	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		-- Write strobes. This signal indicates which byte lanes hold
    		-- valid data. There is one write strobe bit for each eight
    		-- bits of the write data bus.    
		S_AXI_WSTRB	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		-- Write valid. This signal indicates that valid write
    		-- data and strobes are available.
		S_AXI_WVALID	: in std_logic;
		-- Write ready. This signal indicates that the slave
    		-- can accept the write data.
		S_AXI_WREADY	: out std_logic;
		-- Write response. This signal indicates the status
    		-- of the write transaction.
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		-- Write response valid. This signal indicates that the channel
    		-- is signaling a valid write response.
		S_AXI_BVALID	: out std_logic;
		-- Response ready. This signal indicates that the master
    		-- can accept a write response.
		S_AXI_BREADY	: in std_logic;
		-- Read address (issued by master, acceped by Slave)
		S_AXI_ARADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		-- Protection type. This signal indicates the privilege
    		-- and security level of the transaction, and whether the
    		-- transaction is a data access or an instruction access.
		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		-- Read address valid. This signal indicates that the channel
    		-- is signaling valid read address and control information.
		S_AXI_ARVALID	: in std_logic;
		-- Read address ready. This signal indicates that the slave is
    		-- ready to accept an address and associated control signals.
		S_AXI_ARREADY	: out std_logic;
		-- Read data (issued by slave)
		S_AXI_RDATA	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		-- Read response. This signal indicates the status of the
    		-- read transfer.
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		-- Read valid. This signal indicates that the channel is
    		-- signaling the required read data.
		S_AXI_RVALID	: out std_logic;
		-- Read ready. This signal indicates that the master can
    		-- accept the read data and response information.
		S_AXI_RREADY	: in std_logic
	);
end laelaps_four_legs_duplicate_ip_v1_0_S00_AXI;

architecture arch_imp of laelaps_four_legs_duplicate_ip_v1_0_S00_AXI is

	-- AXI4LITE signals
	signal axi_awaddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_awready	: std_logic;
	signal axi_wready	: std_logic;
	signal axi_bresp	: std_logic_vector(1 downto 0);
	signal axi_bvalid	: std_logic;
	signal axi_araddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_arready	: std_logic;
	signal axi_rdata	: std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal axi_rresp	: std_logic_vector(1 downto 0);
	signal axi_rvalid	: std_logic;

	-- Example-specific design signals
	-- local parameter for addressing 32 bit / 64 bit C_S_AXI_DATA_WIDTH
	-- ADDR_LSB is used for addressing 32/64 bit registers/memories
	-- ADDR_LSB = 2 for 32 bits (n downto 2)
	-- ADDR_LSB = 3 for 64 bits (n downto 3)
	constant ADDR_LSB  : integer := (C_S_AXI_DATA_WIDTH/32)+ 1;
	constant OPT_MEM_ADDR_BITS : integer := 4;
	------------------------------------------------
	---- Signals for user logic register space example
    ------------------------------------------------

    --LEG NUMBER 1
     ---------------
     --FOR QEI
     --signals for ENCODER 1 LEG 1
     signal Counts1_1 : STD_LOGIC_VECTOR (bits-1 downto 0);    --Counts of encoder 1 of leg 1
     signal vel_sign1_1 : std_logic;
     signal vel1_1 : std_logic_vector(31 downto 0);            --Velocity of motor 1 of leg 1
             
     --signals for ENCODER 2 LEG 1
     signal Counts2_1 : STD_LOGIC_VECTOR (bits-1 downto 0);    --Counts of encoder 2 of leg 1
     signal vel_sign2_1 : std_logic;
     signal vel2_1 : std_logic_vector(31 downto 0);            --Velocity of motor 2 of leg 1
     
     --FOR PWM
     signal pwm_output1_1 : std_logic_vector(phases-1 downto 0); --PWM signal for motor 1 of leg 1
     signal pwm_output2_1 : std_logic_vector(phases-1 downto 0); --PWM signal for motor 2 of leg 1
     --------------------------------------------------------------------------------------
     
     --------------------------------------------------------------------------------------
     --LEG NUMBER 2
     ---------------
     --FOR QEI
     --signals for ENCODER 1 LEG 2
     signal Counts1_2 : STD_LOGIC_VECTOR (bits-1 downto 0);    --Counts of encoder 1 of leg 2
     signal vel_sign1_2 : std_logic;
     signal vel1_2 : std_logic_vector(31 downto 0);            --Velocity of motor 1 of leg 2
             
     --signals for ENCODER 2 LEG 2
     signal Counts2_2 : STD_LOGIC_VECTOR (bits-1 downto 0);    --Counts of encoder 2 of leg 2
     signal vel_sign2_2 : std_logic;
     signal vel2_2 : std_logic_vector(31 downto 0);            --Velocity of motor 2 of leg 2
     
     --FOR PWM
     signal pwm_output1_2 : std_logic_vector(phases-1 downto 0); --PWM signal for motor 1 of leg 2
     signal pwm_output2_2 : std_logic_vector(phases-1 downto 0); --PWM signal for motor 2 of leg 2
     ----------------------------------------------------------------------------------------------
     --------------------------------------------------------------------------------------
     --LEG NUMBER 3
     ---------------
     --FOR QEI
     --signals for ENCODER 1 LEG 3
     signal Counts1_3 : STD_LOGIC_VECTOR (bits-1 downto 0);    --Counts of encoder 1 of leg 3
     signal vel_sign1_3 : std_logic;
     signal vel1_3 : std_logic_vector(31 downto 0);            --Velocity of motor 1 of leg 3
             
     --signals for ENCODER 2 LEG 3
     signal Counts2_3 : STD_LOGIC_VECTOR (bits-1 downto 0);    --Counts of encoder 2 of leg 3
     signal vel_sign2_3 : std_logic;
     signal vel2_3 : std_logic_vector(31 downto 0);            --Velocity of motor 2 of leg 3
     
     --FOR PWM
     signal pwm_output1_3 : std_logic_vector(phases-1 downto 0); --PWM signal for motor 1 of leg 3
     signal pwm_output2_3 : std_logic_vector(phases-1 downto 0); --PWM signal for motor 2 of leg 3
     ----------------------------------------------------------------------------------------------
     --------------------------------------------------------------------------------------
     --LEG NUMBER 4
     ---------------
     --FOR QEI
     --signals for ENCODER 1 LEG 4
     signal Counts1_4 : STD_LOGIC_VECTOR (bits-1 downto 0);    --Counts of encoder 1 of leg 4
     signal vel_sign1_4 : std_logic;
     signal vel1_4 : std_logic_vector(31 downto 0);            --Velocity of motor 1 of leg 4
             
     --signals for ENCODER 2 LEG 4
     signal Counts2_4 : STD_LOGIC_VECTOR (bits-1 downto 0);    --Counts of encoder 2 of leg 4
     signal vel_sign2_4 : std_logic;
     signal vel2_4 : std_logic_vector(31 downto 0);            --Velocity of motor 2 of leg 4
     
     --FOR PWM
     signal pwm_output1_4 : std_logic_vector(phases-1 downto 0); --PWM signal for motor 1 of leg 4
     signal pwm_output2_4 : std_logic_vector(phases-1 downto 0); --PWM signal for motor 2 of leg 4
     ----------------------------------------------------------------------------------------------
     -- Auxiliary signals
     signal led0_temp0 : std_logic_vector(phases-1 downto 0);
     signal led0_temp1 : std_logic_vector(phases-1 downto 0);
     signal led0_temp2 : std_logic_vector(phases-1 downto 0);
     signal led0_temp3 : std_logic_vector(phases-1 downto 0);
     
     signal led1_temp0 : std_logic;
     signal led1_temp1 : std_logic;
     signal led1_temp2 : std_logic;
     signal led1_temp3 : std_logic;
 
     signal led2_temp0 : std_logic_vector(phases-1 downto 0);
     signal led2_temp1 : std_logic_vector(phases-1 downto 0);
     signal led2_temp2 : std_logic_vector(phases-1 downto 0);
     signal led2_temp3 : std_logic_vector(phases-1 downto 0);
 
     signal led3_temp0 : std_logic;
     signal led3_temp1 : std_logic;
     signal led3_temp2 : std_logic;
     signal led3_temp3 : std_logic;
     
     ----------------------------------------------------------------------------------------------
     --Declaration of components
     component qei
        generic(--these are not the actual values of the generic variables. See Generic Map Lines 486 & 502
            sys_clk         : INTEGER := 100_000_000;           --system clock frequency in Hz
            bits            : INTEGER := 18;                    --number of ratio bits
            ratio_numerator : INTEGER := 98;                    --numerator of the gear ratio of the motor-gearhead
            ratio_divisor   : INTEGER := 1                      --divisor of the gear ratio of the motor-gearhead
             ); 
        Port ( 
            QEA : in STD_LOGIC;                                  --The A signal as generated from the encoder
            Index : in STD_LOGIC;                                --The Index signal as generated from the encoder
            QEB : in STD_LOGIC;                                  --The B signal as generated from the encoder
            Clk : in STD_LOGIC;                                  --The Clock Signal
            Count_out : out STD_LOGIC_VECTOR (bits-1 downto 0);  --The Calculated Position of the Motor in Counts
            vel_sign : out STD_LOGIC;                            --The Calculated Sign of the Motor's Velocity
            velocity : out STD_LOGIC_VECTOR  (31 downto 0)       --The Calculated Value of the Motor's Velocity
            );
     end component;  
     
     component pwm_freq IS
        GENERIC(              --The values defined below will only apply in case the "pwm_freq" entity is used as the top module
                              --Otherwise, if another project utilizes it as a component, then the generic variables will be defined there (See the corresponding "Generic Map")
            sys_clk         : INTEGER := 100_000_000;                             --system's clock frequency in Hz
            pwm_frequency   : INTEGER := 20_000;                                  --PWM switching frequency in Hz
            bits_resolution : INTEGER := 14;                                      --bits of resolution setting the duty cycle
            phases          : INTEGER := 1);                                      --number of output pwms and phases
        PORT(
            clk       : IN  STD_LOGIC;                                            --system clock
            reset     : IN  STD_LOGIC;                                            --asynchronous reset
            ena       : IN  STD_LOGIC;                                            --latches in new duty cycle
            duty      : IN  STD_LOGIC_VECTOR(bits_resolution-1 DOWNTO 0);         --duty cycle
            pwm_out   : OUT STD_LOGIC_VECTOR(phases-1 DOWNTO 0));                 --pwm outputs
     END component; 
     ------------------------------------------------
	--------------------------------------------------
	---- Number of Slave Registers 24
	signal slv_reg0	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg1	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg2	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg3	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg4	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg5	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg6	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg7	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg8	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg9	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg10	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg11	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg12	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg13	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg14	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg15	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg16	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg17	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg18	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg19	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg20	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg21	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg22	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg23	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg_rden	: std_logic;
	signal slv_reg_wren	: std_logic;
	signal reg_data_out	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal byte_index	: integer;
	signal aw_en	: std_logic;

begin
	-- I/O Connections assignments

	S_AXI_AWREADY	<= axi_awready;
	S_AXI_WREADY	<= axi_wready;
	S_AXI_BRESP	<= axi_bresp;
	S_AXI_BVALID	<= axi_bvalid;
	S_AXI_ARREADY	<= axi_arready;
	S_AXI_RDATA	<= axi_rdata;
	S_AXI_RRESP	<= axi_rresp;
	S_AXI_RVALID	<= axi_rvalid;
	-- Implement axi_awready generation
	-- axi_awready is asserted for one S_AXI_ACLK clock cycle when both
	-- S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
	-- de-asserted when reset is low.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awready <= '0';
	      aw_en <= '1';
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1' and aw_en = '1') then
	        -- slave is ready to accept write address when
	        -- there is a valid write address and write data
	        -- on the write address and data bus. This design 
	        -- expects no outstanding transactions. 
	        axi_awready <= '1';
	        elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then
	            aw_en <= '1';
	        	axi_awready <= '0';
	      else
	        axi_awready <= '0';
	      end if;
	    end if;
	  end if;
	end process;

	-- Implement axi_awaddr latching
	-- This process is used to latch the address when both 
	-- S_AXI_AWVALID and S_AXI_WVALID are valid. 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awaddr <= (others => '0');
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1' and aw_en = '1') then
	        -- Write Address latching
	        axi_awaddr <= S_AXI_AWADDR;
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement axi_wready generation
	-- axi_wready is asserted for one S_AXI_ACLK clock cycle when both
	-- S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_wready is 
	-- de-asserted when reset is low. 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_wready <= '0';
	    else
	      if (axi_wready = '0' and S_AXI_WVALID = '1' and S_AXI_AWVALID = '1' and aw_en = '1') then
	          -- slave is ready to accept write data when 
	          -- there is a valid write address and write data
	          -- on the write address and data bus. This design 
	          -- expects no outstanding transactions.           
	          axi_wready <= '1';
	      else
	        axi_wready <= '0';
	      end if;
	    end if;
	  end if;
	end process; 

	-- Implement memory mapped register select and write logic generation
	-- The write data is accepted and written to memory mapped registers when
	-- axi_awready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted. Write strobes are used to
	-- select byte enables of slave registers while writing.
	-- These registers are cleared when reset (active low) is applied.
	-- Slave register write enable is asserted when valid address and data are available
	-- and the slave is ready to accept the write address and write data.
	slv_reg_wren <= axi_wready and S_AXI_WVALID and axi_awready and S_AXI_AWVALID ;

	process (S_AXI_ACLK)
	variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS downto 0); 
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      slv_reg0 <= (others => '0');
	      slv_reg1 <= (others => '0');
	      slv_reg2 <= (others => '0');
	      slv_reg3 <= (others => '0');
	      slv_reg4 <= (others => '0');
	      slv_reg5 <= (others => '0');
	      slv_reg6 <= (others => '0');
	      slv_reg7 <= (others => '0');
	      slv_reg8 <= (others => '0');
	      slv_reg9 <= (others => '0');
	      slv_reg10 <= (others => '0');
	      slv_reg11 <= (others => '0');
	      slv_reg12 <= (others => '0');
	      slv_reg13 <= (others => '0');
	      slv_reg14 <= (others => '0');
	      slv_reg15 <= (others => '0');
	      slv_reg16 <= (others => '0');
	      slv_reg17 <= (others => '0');
	      slv_reg18 <= (others => '0');
	      slv_reg19 <= (others => '0');
	      slv_reg20 <= (others => '0');
	      slv_reg21 <= (others => '0');
	      slv_reg22 <= (others => '0');
	      slv_reg23 <= (others => '0');
	    else
	      loc_addr := axi_awaddr(ADDR_LSB + OPT_MEM_ADDR_BITS downto ADDR_LSB);
	      if (slv_reg_wren = '1') then
	        case loc_addr is
	          when b"00000" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 0
	                slv_reg0(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00001" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 1
	                slv_reg1(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00010" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 2
	                slv_reg2(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00011" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 3
	                slv_reg3(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00100" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 4
	                slv_reg4(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00101" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 5
	                slv_reg5(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00110" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 6
	                slv_reg6(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00111" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 7
	                slv_reg7(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01000" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 8
	                slv_reg8(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01001" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 9
	                slv_reg9(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01010" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 10
	                slv_reg10(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01011" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 11
	                slv_reg11(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01100" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 12
	                slv_reg12(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01101" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 13
	                slv_reg13(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01110" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 14
	                slv_reg14(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01111" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 15
	                slv_reg15(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10000" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 16
	                slv_reg16(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10001" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 17
	                slv_reg17(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10010" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 18
	                slv_reg18(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10011" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 19
	                slv_reg19(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10100" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 20
	                slv_reg20(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10101" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 21
	                slv_reg21(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10110" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 22
	                slv_reg22(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10111" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 23
	                slv_reg23(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when others =>
	            slv_reg0 <= slv_reg0;
	            slv_reg1 <= slv_reg1;
	            slv_reg2 <= slv_reg2;
	            slv_reg3 <= slv_reg3;
	            slv_reg4 <= slv_reg4;
	            slv_reg5 <= slv_reg5;
	            slv_reg6 <= slv_reg6;
	            slv_reg7 <= slv_reg7;
	            slv_reg8 <= slv_reg8;
	            slv_reg9 <= slv_reg9;
	            slv_reg10 <= slv_reg10;
	            slv_reg11 <= slv_reg11;
	            slv_reg12 <= slv_reg12;
	            slv_reg13 <= slv_reg13;
	            slv_reg14 <= slv_reg14;
	            slv_reg15 <= slv_reg15;
	            slv_reg16 <= slv_reg16;
	            slv_reg17 <= slv_reg17;
	            slv_reg18 <= slv_reg18;
	            slv_reg19 <= slv_reg19;
	            slv_reg20 <= slv_reg20;
	            slv_reg21 <= slv_reg21;
	            slv_reg22 <= slv_reg22;
	            slv_reg23 <= slv_reg23;
	        end case;
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement write response logic generation
	-- The write response and response valid signals are asserted by the slave 
	-- when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
	-- This marks the acceptance of address and indicates the status of 
	-- write transaction.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_bvalid  <= '0';
	      axi_bresp   <= "00"; --need to work more on the responses
	    else
	      if (axi_awready = '1' and S_AXI_AWVALID = '1' and axi_wready = '1' and S_AXI_WVALID = '1' and axi_bvalid = '0'  ) then
	        axi_bvalid <= '1';
	        axi_bresp  <= "00"; 
	      elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then   --check if bready is asserted while bvalid is high)
	        axi_bvalid <= '0';                                 -- (there is a possibility that bready is always asserted high)
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement axi_arready generation
	-- axi_arready is asserted for one S_AXI_ACLK clock cycle when
	-- S_AXI_ARVALID is asserted. axi_awready is 
	-- de-asserted when reset (active low) is asserted. 
	-- The read address is also latched when S_AXI_ARVALID is 
	-- asserted. axi_araddr is reset to zero on reset assertion.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_arready <= '0';
	      axi_araddr  <= (others => '1');
	    else
	      if (axi_arready = '0' and S_AXI_ARVALID = '1') then
	        -- indicates that the slave has acceped the valid read address
	        axi_arready <= '1';
	        -- Read Address latching 
	        axi_araddr  <= S_AXI_ARADDR;           
	      else
	        axi_arready <= '0';
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement axi_arvalid generation
	-- axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both 
	-- S_AXI_ARVALID and axi_arready are asserted. The slave registers 
	-- data are available on the axi_rdata bus at this instance. The 
	-- assertion of axi_rvalid marks the validity of read data on the 
	-- bus and axi_rresp indicates the status of read transaction.axi_rvalid 
	-- is deasserted on reset (active low). axi_rresp and axi_rdata are 
	-- cleared to zero on reset (active low).  
	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then
	    if S_AXI_ARESETN = '0' then
	      axi_rvalid <= '0';
	      axi_rresp  <= "00";
	    else
	      if (axi_arready = '1' and S_AXI_ARVALID = '1' and axi_rvalid = '0') then
	        -- Valid read data is available at the read data bus
	        axi_rvalid <= '1';
	        axi_rresp  <= "00"; -- 'OKAY' response
	      elsif (axi_rvalid = '1' and S_AXI_RREADY = '1') then
	        -- Read data is accepted by the master
	        axi_rvalid <= '0';
	      end if;            
	    end if;
	  end if;
	end process;

	-- Implement memory mapped register select and read logic generation
	-- Slave register read enable is asserted when valid address is available
	-- and the slave is ready to accept the read address.
	slv_reg_rden <= axi_arready and S_AXI_ARVALID and (not axi_rvalid) ;

	process (Counts1_1, vel_sign1_1, vel1_1, slv_reg2, Counts2_1, vel_sign2_1, vel2_1, slv_reg5, Counts1_2, vel_sign1_2, vel1_2, slv_reg8, Counts2_2, vel_sign2_2, vel2_2, slv_reg11, Counts1_3, vel_sign1_3, vel1_3, slv_reg14, Counts2_3, vel_sign2_3, vel2_3, slv_reg17, Counts1_4, vel_sign1_4, vel1_4, slv_reg20, Counts2_4, vel_sign2_4, vel2_4, slv_reg23, axi_araddr, S_AXI_ARESETN, slv_reg_rden)
	variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS downto 0);
	begin
        -- Address decoding for reading registers
        loc_addr := axi_araddr(ADDR_LSB + OPT_MEM_ADDR_BITS downto ADDR_LSB);
        case loc_addr is
          when b"00000" =>
--            reg_data_out <= slv_reg0;
            reg_data_out(31 downto bits+1) <= (others => '0');
            reg_data_out(bits) <= vel_sign1_1;                  --Send the Sign of velocity for motor 1 leg 1
            reg_data_out(bits-1 downto 0 ) <= Counts1_1;        --Send the Counter of QEI for encoder 1 leg 1
          when b"00001" =>
--            reg_data_out <= slv_reg1;
            reg_data_out(31 downto 0 ) <= vel1_1;               --Send the Velocity of motor 1 leg 1          
          when b"00010" =>
            reg_data_out <= slv_reg2;                           --Read the register relevant with the PWM of motor 1 leg 1
          when b"00011" =>
--            reg_data_out <= slv_reg3;
            reg_data_out(31 downto bits+1) <= (others => '0');
            reg_data_out(bits) <= vel_sign2_1;                  --Send the Sign of velocity for motor 2 leg 1
            reg_data_out(bits-1 downto 0 ) <= Counts2_1;        --Send the Counter of QEI for encoder 2 leg 1
          when b"00100" =>
--            reg_data_out <= slv_reg4;
            reg_data_out(31 downto 0 ) <= vel2_1;               --Send the Velocity of motor 2 leg 1
          when b"00101" =>
            reg_data_out <= slv_reg5;                           --Read the egister relevant with the PWM of motor 2 leg 1
          when b"00110" =>
--            reg_data_out <= slv_reg6;
            reg_data_out(31 downto bits+1) <= (others => '0');
            reg_data_out(bits) <= vel_sign1_2;                  --Send the Sign of velocity for motor 1 leg 2
            reg_data_out(bits-1 downto 0 ) <= Counts1_2;        --Send the Counter of QEI for encoder 1 leg 2
          when b"00111" =>
--            reg_data_out <= slv_reg7;
            reg_data_out(31 downto 0 ) <= vel1_2;               --Send the Velocity of motor 1 leg 2
          when b"01000" =>
            reg_data_out <= slv_reg8;                           --Read the register relevant with the PWM of motor 1 leg 2
          when b"01001" =>
--            reg_data_out <= slv_reg9;
            reg_data_out(31 downto bits+1) <= (others => '0');
            reg_data_out(bits) <= vel_sign2_2;                  --Send the Sign of velocity for motor 2 leg 2
            reg_data_out(bits-1 downto 0 ) <= Counts2_2;        --Send the Counter of QEI for encoder 2 leg 2
          when b"01010" =>
--            reg_data_out <= slv_reg10;
            reg_data_out(31 downto 0 ) <= vel2_2;               --Send the Velocity of motor 2 leg 2
          when b"01011" =>
            reg_data_out <= slv_reg11;                          --Read the register relevant with the PWM of motor 2 leg 2
          when b"01100" =>
--            reg_data_out <= slv_reg12;
            reg_data_out(31 downto bits+1) <= (others => '0');
            reg_data_out(bits) <= vel_sign1_3;                  --Send the Sign of velocity for motor 1 leg 3
            reg_data_out(bits-1 downto 0 ) <= Counts1_3;        --Send the Counter of QEI for encoder 1 leg 3
          when b"01101" =>
--            reg_data_out <= slv_reg13;
            reg_data_out(31 downto 0 ) <= vel1_3;               --Send the Velocity of motor 1 leg 3
          when b"01110" =>
            reg_data_out <= slv_reg14;                          --Read the register relevant with the PWM of motor 1 leg 3               
          when b"01111" =>
--            reg_data_out <= slv_reg15;
            reg_data_out(31 downto bits+1) <= (others => '0');
            reg_data_out(bits) <= vel_sign2_3;                  --Send the Sign of velocity for motor 2 leg 3
            reg_data_out(bits-1 downto 0 ) <= Counts2_3;        --Send the Counter of QEI for encoder 2 leg 3
          when b"10000" =>
--            reg_data_out <= slv_reg16;
            reg_data_out(31 downto 0 ) <= vel2_3;               --Send the Velocity of motor 2 leg 3
          when b"10001" =>
            reg_data_out <= slv_reg17;                          --Read the register relevant with the PWM of motor 2 leg 3
          when b"10010" =>
--            reg_data_out <= slv_reg18;
            reg_data_out(31 downto bits+1) <= (others => '0');
            reg_data_out(bits) <= vel_sign1_4;                  --Send the Sign of velocity for motor 1 leg 4
            reg_data_out(bits-1 downto 0 ) <= Counts1_4;        --Send the Counter of QEI for encoder 1 leg 4
          when b"10011" =>
--            reg_data_out <= slv_reg19;
            reg_data_out(31 downto 0 ) <= vel1_4;               --Send the Velocity of motor 1 leg 4
          when b"10100" =>
            reg_data_out <= slv_reg20;                          --Read the register relevant with the PWM of motor 1 leg 4
          when b"10101" =>
--            reg_data_out <= slv_reg21;
            reg_data_out(31 downto bits+1) <= (others => '0');
            reg_data_out(bits) <= vel_sign2_4;                  --Send the Sign of velocity for motor 2 leg 4
            reg_data_out(bits-1 downto 0 ) <= Counts2_4;        --Send the Counter of QEI for encoder 2 leg 4
          when b"10110" =>
--            reg_data_out <= slv_reg22;
            reg_data_out(31 downto 0 ) <= vel2_4;               --Send the Velocity of motor 2 leg 4
          when b"10111" =>
            reg_data_out <= slv_reg23;                          --Read the register relevant with the PWM of motor 2 leg 4
          when others =>
            reg_data_out  <= (others => '0');
        end case;
    end process; 

	-- Output register or memory read data
	process( S_AXI_ACLK ) is
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	      axi_rdata  <= (others => '0');
	    else
	      if (slv_reg_rden = '1') then
	        -- When there is a valid read address (S_AXI_ARVALID) with 
	        -- acceptance of read address by the slave (axi_arready), 
	        -- output the read dada 
	        -- Read address mux
	          axi_rdata <= reg_data_out;     -- register read data
	      end if;   
	    end if;
	  end if;
	end process;


	-- Add user logic here
--QEIs start here
    cl1: qei                                                    --QEI for motor-encoder 1 leg 1
        generic map(sys_clk => sys_clk, 
                    bits => bits,
                    ratio_numerator => hip_ratio_numerator,
                    ratio_divisor => hip_ratio_divisor
                    )
        port map(
            QEA => jb_p0,
            Index => '0',
            QEB => jb_n0,
            Clk => S_AXI_ACLK,
            Count_out => Counts1_1,
            vel_sign => vel_sign1_1,
            velocity => vel1_1
        );
                        
    cl2: qei                                                    --QEI for motor-encoder 2 leg 1         
        generic map(sys_clk => sys_clk, 
                    bits => bits,
                    ratio_numerator => knee_ratio_numerator,
                    ratio_divisor => knee_ratio_divisor
                    )
        port map(
            QEA => jb_p1,
            Index => '0',
            QEB => jb_n1,
            Clk => S_AXI_ACLK,
            Count_out => Counts2_1,
            vel_sign => vel_sign2_1,
            velocity => vel2_1
        ); 
    
    cl3: qei                                                    --QEI for motor-encoder 1 leg 2
        generic map(sys_clk => sys_clk, 
                    bits => bits,
                    ratio_numerator => hip_ratio_numerator,
                    ratio_divisor => hip_ratio_divisor
                    )
        port map(
            QEA => jc_p0,
            Index => '0',
            QEB => jc_n0,
            Clk => S_AXI_ACLK,
            Count_out => Counts1_2,
            vel_sign => vel_sign1_2,
            velocity => vel1_2
        );
                        
    cl4: qei                                                    --QEI for motor-encoder 2 leg 2         
        generic map(sys_clk => sys_clk, 
                    bits => bits,
                    ratio_numerator => knee_ratio_numerator,
                    ratio_divisor => knee_ratio_divisor
                    )
        port map(
            QEA => jc_p1,
            Index => '0',
            QEB => jc_n1,
            Clk => S_AXI_ACLK,
            Count_out => Counts2_2,
            vel_sign => vel_sign2_2,
            velocity => vel2_2
        ); 
            
    cl5: qei                                                    --QEI for motor-encoder 1 leg 3
        generic map(sys_clk => sys_clk, 
                    bits => bits,
                    ratio_numerator => hip_ratio_numerator,
                    ratio_divisor => hip_ratio_divisor
                    )
        port map(
            QEA => jd_p0,
            Index => '0',
            QEB => jd_n0,
            Clk => S_AXI_ACLK,
            Count_out => Counts1_3,
            vel_sign => vel_sign1_3,
            velocity => vel1_3
        );
                        
    cl6: qei                                                    --QEI for motor-encoder 2 leg 3         
        generic map(sys_clk => sys_clk, 
                    bits => bits,
                    ratio_numerator => knee_ratio_numerator,
                    ratio_divisor => knee_ratio_divisor
                    )
        port map(
            QEA => jd_p1,
            Index => '0',
            QEB => jd_n1,
            Clk => S_AXI_ACLK,
            Count_out => Counts2_3,
            vel_sign => vel_sign2_3,
            velocity => vel2_3
        ); 
    
    cl7: qei                                                    --QEI for motor-encoder 1 leg 4
        generic map(sys_clk => sys_clk, 
                    bits => bits,
                    ratio_numerator => hip_ratio_numerator,
                    ratio_divisor => hip_ratio_divisor
                    )
        port map(
            QEA => je_p0,
            Index => '0',
            QEB => je_n0,
            Clk => S_AXI_ACLK,
            Count_out => Counts1_4,
            vel_sign => vel_sign1_4,
            velocity => vel1_4
        );
                        
    cl8: qei                                                    --QEI for motor-encoder 2 leg 4         
        generic map(sys_clk => sys_clk, 
                    bits => bits,
                    ratio_numerator => knee_ratio_numerator,
                    ratio_divisor => knee_ratio_divisor
                    )
        port map(
            QEA => je_p1,
            Index => '0',
            QEB => je_n1,
            Clk => S_AXI_ACLK,
            Count_out => Counts2_4,
            vel_sign => vel_sign2_4,
            velocity => vel2_4
        );
    --QEIs end here
    
    --PWMs start here
    
    --LEG NUMBER 1
    pwm_freq_1 : pwm_freq                                       --PWM for motor 1 leg 1
        generic map (sys_clk => sys_clk,                        --system clock frequency in Hz
              pwm_frequency => pwm_frequency,                   --PWM switching frequency in Hz
              bits_resolution => bits_resolution,               --bits of resolution setting the duty cycle
              phases          => phases                         --number of output pwms and phases
            )
        port map(
            clk => S_AXI_ACLK,                                  --system clock
            reset  => slv_reg2(0),                              --Asynchronous reset of duty cycle for Motor 1 Leg 1
            ena  => slv_reg2(1),                                --Latches in new duty cycle for Motor 1 Leg 1
            duty => slv_reg2(bits_resolution-1+3 downto 3),     --Duty cycle for Motor 1 Leg 1
            pwm_out  => pwm_output1_1                           --Pwm output for Motor 1 Leg 1
        );
        
        jb_p2 <= slv_reg2(2);                                   --Direction Signal for Motor 1 Leg 1
        jb_n2 <= pwm_output1_1(0);                              --PWM Signal for Motor 1 Leg 1
                  
    pwm_freq_2 : pwm_freq                                       --PWM for motor 2 leg 1
        generic map (sys_clk => sys_clk,                        --system clock frequency in Hz
              pwm_frequency => pwm_frequency,                   --PWM switching frequency in Hz
              bits_resolution => bits_resolution,               --bits of resolution setting the duty cycle
              phases          => phases                         --number of output pwms and phases
        )
        port map(
                clk => S_AXI_ACLK,                              --system clock
                reset  => slv_reg5(0),                          --Asynchronous reset of duty cycle for Motor 2 Leg 1
                ena  => slv_reg5(1),                            --Latches in new duty cycle for Motor 2 Leg 1
                duty => slv_reg5(bits_resolution-1+3 downto 3), --Duty cycle for Motor 2 Leg 1
                pwm_out  => pwm_output2_1                       --Pwm output for Motor 2 Leg 1
            );
        
        jb_p3 <= slv_reg5(2);                                   --Direction Signal for Motor 2 Leg 1
        jb_n3 <= pwm_output2_1(0);                              --PWM Signal for Motor 2 Leg 1
    
    --LEG NUMBER 2
    pwm_freq_3 : pwm_freq                                       --PWM for motor 1 leg 2
        generic map (sys_clk => sys_clk,                        --system clock frequency in Hz
              pwm_frequency => pwm_frequency,                   --PWM switching frequency in Hz
              bits_resolution => bits_resolution,               --bits of resolution setting the duty cycle
              phases          => phases                         --number of output pwms and phases
            )
        port map(
            clk => S_AXI_ACLK,                                  --system clock
            reset  => slv_reg8(0),                              --Asynchronous reset of duty cycle for Motor 1 Leg 2
            ena  => slv_reg8(1),                                --Latches in new duty cycle for Motor 1 Leg 2
            duty => slv_reg8(bits_resolution-1+3 downto 3),     --Duty cycle for Motor 1 Leg 2
            pwm_out  => pwm_output1_2                           --Pwm output for Motor 1 Leg 2
        );
        
        jc_p2 <= slv_reg8(2);                                   --Direction Signal for Motor 1 Leg 2
        jc_n2 <= pwm_output1_2(0);                              --PWM Signal for Motor 1 Leg 2
                  
    pwm_freq_4 : pwm_freq                                       --PWM for motor 2 leg 2
        generic map (sys_clk => sys_clk,                        --system clock frequency in Hz
              pwm_frequency => pwm_frequency,                   --PWM switching frequency in Hz
              bits_resolution => bits_resolution,               --bits of resolution setting the duty cycle
              phases          => phases                         --number of output pwms and phases
        )
        port map(
                clk => S_AXI_ACLK,                              --system clock
                reset  => slv_reg11(0),                         --Asynchronous reset of duty cycle for Motor 2 Leg 2
                ena  => slv_reg11(1),                           --Latches in new duty cycle for Motor 2 Leg 2
                duty => slv_reg11(bits_resolution-1+3 downto 3),--Duty cycle for Motor 2 Leg 2
                pwm_out  => pwm_output2_2                       --Pwm output for Motor 2 Leg 2
            );
        
        jc_p3 <= slv_reg11(2);                                  --Direction Signal for Motor 2 Leg 2
        jc_n3 <= pwm_output2_2(0);                              --PWM Signal for Motor 2 Leg 2
    ---
    --LEG NUMBER 3
    pwm_freq_5 : pwm_freq                                       --PWM for motor 1 leg 3
        generic map (sys_clk => sys_clk,                        --system clock frequency in Hz
              pwm_frequency => pwm_frequency,                   --PWM switching frequency in Hz
              bits_resolution => bits_resolution,               --bits of resolution setting the duty cycle
              phases          => phases                         --number of output pwms and phases
            )
        port map(
            clk => S_AXI_ACLK,                                  --system clock
            reset  => slv_reg14(0),                             --Asynchronous reset of duty cycle for Motor 1 Leg 3
            ena  => slv_reg14(1),                               --Latches in new duty cycle for Motor 1 Leg 3
            duty => slv_reg14(bits_resolution-1+3 downto 3),    --Duty cycle for Motor 1 Leg 3
            pwm_out  => pwm_output1_3                           --Pwm output for Motor 1 Leg 3
        );
        
        jd_p2 <= slv_reg14(2);                                  --Direction Signal for Motor 1 Leg 3
        jd_n2 <= pwm_output1_3(0);                              --PWM Signal for Motor 1 Leg 3
                  
    pwm_freq_6 : pwm_freq                                       --PWM for motor 2 leg 3
        generic map (sys_clk => sys_clk,                        --system clock frequency in Hz
              pwm_frequency => pwm_frequency,                   --PWM switching frequency in Hz
              bits_resolution => bits_resolution,               --bits of resolution setting the duty cycle
              phases          => phases                         --number of output pwms and phases
        )
        port map(
                clk => S_AXI_ACLK,                              --system clock
                reset  => slv_reg17(0),                         --Asynchronous reset of duty cycle for Motor 2 Leg 3
                ena  => slv_reg17(1),                           --Latches in new duty cycle for Motor 2 Leg 3
                duty => slv_reg17(bits_resolution-1+3 downto 3),--Duty cycle for Motor 2 Leg 3
                pwm_out  => pwm_output2_3                       --Pwm output for Motor 2 Leg 3
            );
        
        jd_p3 <= slv_reg17(2);                                   --Direction Signal for Motor 2 Leg 3
        jd_n3 <= pwm_output2_3(0);                              --PWM Signal for Motor 2 Leg 3
    
    --LEG NUMBER 4
    pwm_freq_7 : pwm_freq                                       --PWM for motor 1 leg 4
        generic map (sys_clk => sys_clk,                        --system clock frequency in Hz
              pwm_frequency => pwm_frequency,                   --PWM switching frequency in Hz
              bits_resolution => bits_resolution,               --bits of resolution setting the duty cycle
              phases          => phases                         --number of output pwms and phases
            )
        port map(
            clk => S_AXI_ACLK,                                  --system clock
            reset  => slv_reg20(0),                              --Asynchronous reset of duty cycle for Motor 1 Leg 4
            ena  => slv_reg20(1),                                --Latches in new duty cycle for Motor 1 Leg 4
            duty => slv_reg20(bits_resolution-1+3 downto 3),     --Duty cycle for Motor 1 Leg 4
            pwm_out  => pwm_output1_4                           --Pwm output for Motor 1 Leg 4
        );
        
        je_p2 <= slv_reg20(2);                                   --Direction Signal for Motor 1 Leg 4
        je_n2 <= pwm_output1_4(0);                              --PWM Signal for Motor 1 Leg 4
                  
    pwm_freq_8 : pwm_freq                                       --PWM for motor 2 leg 4
        generic map (sys_clk => sys_clk,                        --system clock frequency in Hz
              pwm_frequency => pwm_frequency,                   --PWM switching frequency in Hz
              bits_resolution => bits_resolution,               --bits of resolution setting the duty cycle
              phases          => phases                         --number of output pwms and phases
        )
        port map(
                clk => S_AXI_ACLK,                              --system clock
                reset  => slv_reg23(0),                         --Asynchronous reset of duty cycle for Motor 2 Leg 4
                ena  => slv_reg23(1),                           --Latches in new duty cycle for Motor 2 Leg 4
                duty => slv_reg23(bits_resolution-1+3 downto 3),--Duty cycle for Motor 2 Leg 4
                pwm_out  => pwm_output2_4                       --Pwm output for Motor 2 Leg 4
            );
        
        je_p3 <= slv_reg23(2);                                  --Direction Signal for Motor 2 Leg 4
        je_n3 <= pwm_output2_4(0);                              --PWM Signal for Motor 2 Leg 4
        
    --PWMs end here
        led0_temp0 <= pwm_output1_1 and sw(phases-1 downto 0);
        led0_temp1 <= pwm_output1_2 and sw(phases downto 1);
        led0_temp2 <= pwm_output1_3 and sw(phases+1 downto 2);
        led0_temp3 <= pwm_output1_4 and sw(phases+2 downto 3);   
       
        led1_temp0 <= slv_reg2(2) and sw(0);
        led1_temp1 <= slv_reg8(2) and sw(1);
        led1_temp2 <= slv_reg2(2) and sw(2);
        led1_temp3 <= slv_reg8(2) and sw(3);
        
        led2_temp0 <= pwm_output2_1 and sw(phases-1 downto 0);
        led2_temp1 <= pwm_output2_2 and sw(phases downto 1);
        led2_temp2 <= pwm_output2_3 and sw(phases+1 downto 2);
        led2_temp3 <= pwm_output2_4 and sw(phases+2 downto 3);
            
        led3_temp0 <= slv_reg5(2) and sw(0);
        led3_temp1 <= slv_reg11(2) and sw(1);
        led3_temp2 <= slv_reg5(2) and sw(2);
        led3_temp3 <= slv_reg11(2) and sw(3);
        
        led(phases-1 downto 0) <= led0_temp0 or led0_temp1 or led0_temp2 or led0_temp3;      --PWM Signal for Motor 1 of either Leg 1,2,3 or 4 to the first LED of ZYBO
        led(1) <= led1_temp0 or led1_temp1 or led1_temp2 or led1_temp3;                      --Direction Signal for Motor 1 of either Leg 1,2,3 or 4 to the second LED of ZYBO
        led(phases+1 downto 2) <= led2_temp0 or led2_temp1 or led2_temp2 or led2_temp3;      --PWM Signal for Motor 1 of either Leg 1,2,3 or 4 to the third LED of ZYBO
        led(3) <= led3_temp0 or led3_temp1 or led3_temp2 or led3_temp3;                      --Direction Signal for Motor 1 of either Leg 1,2,3 or 4 to the fourth LED of ZYBO
        -- User logic ends

end arch_imp;
